----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08/11/2024 05:46:15 PM
-- Design Name: 
-- Module Name: apply_gaussian_top_simple_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_arith.all;
-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity apply_gaussian_top_simple_tb is
--  Port ( );
end apply_gaussian_top_simple_tb;

architecture Behavioral of apply_gaussian_top_simple_tb is
    constant DRAM_DATA_WIDTH: positive := 8;
 --   constant DRAM_ADDR_WIDTH: positive := 22;
    constant DRAM_SIZE: positive := 6480;
    
    type ram_type is array(0 to DRAM_SIZE-1) of std_logic_vector(DRAM_DATA_WIDTH - 1 downto 0);
    constant DRAM_CONTENT: ram_type := (
B"10001101", B"10000111", B"10000100", B"10001110", B"10100000", B"10101101", B"10110000", B"10101110", B"10011011", B"10010010", B"10001110", B"10001101", B"10001100", B"10001110", B"10010010", B"10010001", B"10010000", B"10001100", B"10001101", B"10001110", B"10001110", B"10001101", B"10010000", B"10011001", B"10100011", B"10101110", B"10110111", B"10110111", B"10101000", B"10010100", B"10001011", B"10001100", B"10001010", B"10000110", B"10000011", B"10000000", B"01111111", B"01111101", B"01111001", B"01111000", B"01111000", B"01111001", B"01111100", B"01111110", B"01111110", B"01111100", B"01111001", B"01111001", B"01111001", B"01111010", B"01111011", B"01111010", B"01111010", B"01111010", B"01111010", B"01111001", B"01111001", B"01111001", B"01111000", B"01111000", B"01110111", B"01110111", B"01110111", B"01110111", B"01111000", B"01111000", B"01110111", B"01110011", B"01110010", B"01110001", B"01110000", B"01110000", B"01101110", B"01101110", B"01101101", B"01101101", B"01101100", B"01101011", B"01101011", B"01101011", B"01101101", B"01101001", B"01101100", B"01101010", B"01110011", B"01110011", B"01001111", B"01000011", B"01011110", B"01101010", B"01101010", B"01101010", B"01110000", B"01110010", B"01101011", B"01110000", B"01110001", B"01111001", B"01110101", B"01110101", B"01110001", B"01110001", B"01111010", B"01110010", B"01110010", B"01100100", B"00110100", B"00100110", B"00110110", B"00111101", B"01000010", B"00111110", B"00111100", B"00111101", B"00111110", B"00111110", B"00111110", B"00111110", B"00111110", B"00111110", B"00111110", B"01000000", B"00111111", B"00110111", B"00101011", B"00100011", B"00100011", B"00100100", B"00100100", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100010", B"00100000", B"00100111", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", 
B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100101", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100111", B"01100111", B"01101000", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", 
B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101010", B"01101010", B"01101011", B"01101011", B"01101100", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101001", B"01101000", B"01101010", B"01101001", B"01100001", B"01011010", B"01100001", B"01110000", B"10011000", B"10010110", B"10010001", B"10001111", B"10010010", B"10010101", B"10011000", B"10010110", B"10010011", B"10010110", B"10011011", B"10011011", B"10011001", B"10011000", B"10011001", B"10011011", B"10011100", B"10011010", B"10011010", B"10011001", B"10011000", B"10010110", B"10010101", B"10010101", B"10010100", B"10010100", B"10010101", B"10010110", B"10011001", B"10011010", B"10011010", B"10011010", B"10011000", B"10010110", B"10010101", B"10010101", B"10010101", B"10010101", B"10010101", B"10010101", B"10010110", B"10010110", B"10011000", B"10011000", B"10011000", B"10011001", B"10011001", B"10011010", B"10011001", B"10010110", B"10010101", B"10010101", B"10010101", B"10010101", B"10010101", B"10010100", B"10010010", B"10001101", B"10001011", B"10001100", B"10001100", B"10001010", B"10000011", B"01111001", B"01101000", B"01011110", B"01101001", B"10000000", B"10001100", B"10000001", B"01110010", B"01101111", B"01111010", B"01111100", B"01111111", B"10000011", B"10000110", B"10001011", B"10001100", B"10001101", B"10001110", B"10001101", B"10001101", B"10001100", B"10001100", B"10001100", B"10001100", B"10001110", B"10011111", B"01111000", B"01010101", B"01001010", B"01001010", B"01001101", B"01010001", B"01010010", B"01001100", B"01110100", B"10010010", B"10010000", B"10001011", B"10010010", B"10010100", B"10001110", B"10000000", B"10000011", B"10001110", B"10001111", B"10001111", B"01101000", B"00111010", B"00111000", B"00110000", B"00100011", B"00011001", B"00100100", B"00110011", B"00101110", B"00110011", B"00110001", B"00111101", B"01000101", B"01001100", B"01010001", B"01010110", B"01011100", B"01101010", B"01111110", B"10000111", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001010", B"10001010", B"10001010", B"10000111", B"10000110", B"10000111", B"10001010", B"10001011", B"10001010", B"10001000", B"10000111", B"10000111", B"10001000", B"10000111", B"10000110", 
B"10000101", B"10000110", B"10001000", B"10001001", B"10001001", B"10001010", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001110", B"10010000", B"10001100", B"01111110", B"01100110", B"01100111", B"01111111", B"10001110", B"10001011", B"10000111", B"10000111", B"10001001", B"10001010", B"10001100", B"10001100", B"10001010", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001010", B"10001100", B"10000011", B"01101011", B"01011011", B"01101001", B"10000011", B"01110110", B"01110011", B"01110001", B"01110010", B"01110001", B"01110000", B"01110001", B"01110001", B"01101000", B"01100000", B"01100100", B"01110110", B"10000001", B"01111111", B"01111010", B"01111001", B"01111010", B"01111010", B"01111100", B"01111101", B"01111101", B"01111110", B"01111110", B"01111110", B"01111110", B"01111111", B"01111111", B"10000000", B"10000000", B"01111110", B"01111101", B"01111110", B"01111000", B"01110001", B"01101110", B"01101011", B"01101011", B"01101001", B"01101010", B"01101001", B"01101000", B"01101000", B"01101010", B"01101100", B"01101111", B"01110001", B"01101100", B"01100101", B"10000110", 
B"10000010", B"10000011", B"10010011", B"10101010", B"10110101", B"10101011", B"10100000", B"10010011", B"10001110", B"10001100", B"10001010", B"10001100", B"10010000", B"10010001", B"10010001", B"10010000", B"10001110", B"10001101", B"10001101", B"10001101", B"10010000", B"10010111", B"10011111", B"10110001", B"10111000", B"11000000", B"10111111", B"10101110", B"10010111", B"10001011", B"10001011", B"10000110", B"10000100", B"10000010", B"10000000", B"01111101", B"01111011", B"01111000", B"01110111", B"01111000", B"01111001", B"01111100", B"01111101", B"01111101", B"01111100", B"01111001", B"01111001", B"01111001", B"01111010", B"01111011", B"01111011", B"01111010", B"01111010", B"01111010", B"01111001", B"01111001", B"01111001", B"01111000", B"01111000", B"01110111", B"01110111", B"01110111", B"01110111", B"01110101", B"01110101", B"01110100", B"01110011", B"01110010", B"01110001", B"01110000", B"01110000", B"01101110", B"01101110", B"01101110", B"01101101", B"01101100", B"01101011", B"01101011", B"01101011", B"01101100", B"01101001", B"01101100", B"01101010", B"01110010", B"01101110", B"01001001", B"01000101", B"01100010", B"01101100", B"01101011", B"01101001", B"01101100", B"01110000", B"01101101", B"01110011", B"01101101", B"01110011", B"01110010", B"01110011", B"01110001", B"01110010", B"01111010", B"01110110", B"01110011", B"01100000", B"00110110", B"00101000", B"00110110", B"00111101", B"00111111", B"00111100", B"00111011", B"00111011", B"00111100", B"00111100", B"00111100", B"00111100", B"00111100", B"00111100", B"00111101", B"00111111", B"00111110", B"00110110", B"00101010", B"00100011", B"00100010", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100010", B"00100000", B"00100111", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", 
B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100101", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100111", B"01100111", B"01101000", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01101000", B"01101000", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", 
B"01101001", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101001", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101000", B"01101010", B"01101001", B"01100001", B"01011010", B"01100001", B"01110000", B"10000110", B"10001100", B"10001101", B"10001100", B"10001000", B"10001011", B"10010011", B"10011001", B"10011000", B"10010110", B"10011001", B"10011000", B"10010101", B"10010011", B"10010101", B"10011000", B"10011000", B"10010110", B"10010110", B"10010110", B"10010101", B"10010101", B"10010100", B"10010011", B"10010011", B"10010011", B"10010011", B"10010101", B"10010110", B"10011000", B"10011000", B"10011000", B"10010110", B"10010101", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010101", B"10010101", B"10010101", B"10010110", B"10010110", B"10010110", B"10010110", B"10010110", B"10010110", B"10010110", B"10010101", B"10010100", B"10010100", B"10010011", B"10010011", B"10010010", B"10001111", B"10001010", B"10001010", B"10001110", B"10010001", B"10010001", B"10000111", B"01111001", B"01101100", B"01011011", B"01100000", B"01111001", B"10010001", B"10010001", B"01111111", B"01110101", B"01110010", B"01100011", B"01100100", B"01100101", B"01100111", B"01101000", B"01101001", B"01101011", B"01101110", B"01110010", B"01110011", B"01110101", B"01110101", B"01110101", B"01110011", B"01110100", B"01110111", B"01110111", B"01100100", B"01010001", B"01001110", B"01010000", B"01001110", B"01001001", B"01000110", B"00111111", B"01101101", B"10001100", B"10001110", B"10001100", B"10010010", B"10010100", B"10001101", B"10011010", B"10011011", B"10011100", B"10001110", B"10000110", B"01100111", B"00111100", B"00101100", B"00011101", B"00011011", B"00011011", B"00100010", B"00100101", B"00011100", B"00101100", B"00111000", B"01001110", B"01001111", B"01010001", B"01011011", B"01011110", B"01100010", B"01110011", B"10000111", B"10010001", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001011", B"10001011", B"10001010", B"10001000", B"10001000", B"10001011", B"10001100", B"10001101", B"10001011", B"10001000", B"10000111", B"10000111", B"10001000", B"10000111", B"10000100", 
B"10000100", B"10000110", B"10001000", B"10001001", B"10001001", B"10001010", B"10001010", B"10001010", B"10001010", B"10001011", B"10001011", B"10001011", B"10001011", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001101", B"10001110", B"10001011", B"01111110", B"01100110", B"01100111", B"01111111", B"10001110", B"10001011", B"10000111", B"10000111", B"10001001", B"10001010", B"10001100", B"10001100", B"10001010", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001010", B"10001100", B"10000011", B"01101011", B"01011011", B"01101001", B"10000011", B"01110110", B"01110010", B"01110001", B"01110001", B"01110001", B"01110000", B"01110001", B"01110001", B"01101000", B"01100000", B"01100100", B"01110110", B"10000000", B"01111111", B"01111001", B"01111000", B"01111001", B"01111010", B"01111010", B"01111100", B"01111100", B"01111101", B"01111101", B"01111101", B"01111101", B"01111101", B"01111101", B"01111110", B"01111101", B"01111010", B"01111001", B"01111010", B"01110010", B"01101110", B"01101001", B"01101000", B"01100111", B"01101000", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101011", B"01101100", B"01101000", B"01100011", B"10000010", 
B"10000100", B"10001110", B"10100000", B"10110000", B"10110001", B"10100010", B"10010100", B"10010010", B"10001110", B"10001011", B"10001011", B"10001101", B"10001101", B"10001101", B"10010000", B"10010010", B"10010001", B"10001110", B"10001100", B"10001110", B"10010111", B"10011111", B"10100111", B"10111011", B"10111110", B"11000110", B"11000101", B"10110001", B"10010101", B"10000110", B"10000111", B"10000101", B"10000011", B"10000010", B"01111111", B"01111011", B"01111000", B"01110111", B"01110101", B"01110111", B"01111001", B"01111100", B"01111010", B"01111010", B"01111100", B"01111010", B"01111010", B"01111011", B"01111011", B"01111100", B"01111011", B"01111010", B"01111010", B"01111010", B"01111001", B"01111001", B"01111001", B"01111001", B"01111000", B"01111000", B"01110111", B"01110101", B"01110101", B"01110101", B"01110100", B"01110100", B"01110011", B"01110010", B"01110001", B"01110000", B"01110000", B"01110000", B"01101101", B"01101101", B"01101100", B"01101100", B"01101011", B"01101010", B"01101011", B"01101010", B"01101010", B"01101100", B"01101011", B"01110001", B"01100110", B"01000001", B"01000111", B"01100111", B"01101110", B"01101011", B"01101001", B"01101010", B"01101101", B"01110001", B"01110111", B"01101011", B"01101111", B"01101110", B"01110000", B"01101110", B"01110000", B"01110100", B"01111000", B"01110000", B"01010110", B"00110101", B"00101101", B"00110110", B"00111110", B"00111111", B"00111110", B"00111101", B"00111101", B"00111101", B"00111100", B"00111100", B"00111100", B"00111100", B"00111100", B"00111100", B"00111101", B"00111011", B"00110101", B"00101010", B"00100011", B"00100010", B"00100010", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100010", B"00100000", B"00100111", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", 
B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100101", B"01100101", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01100101", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101010", B"01101010", B"01101010", 
B"01101001", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01101000", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101000", B"01100111", B"01101001", B"01101000", B"01100000", B"01011001", B"01100000", B"01101010", B"01100011", B"01101011", B"01110101", B"01110101", B"01110000", B"01110010", B"10000000", B"10001100", B"10010110", B"10011100", B"10011111", B"10011011", B"10010110", B"10010100", B"10010100", B"10010101", B"10010101", B"10010110", B"10010110", B"10010110", B"10011000", B"10011000", B"10011000", B"10011000", B"10010110", B"10010101", B"10010101", B"10010110", B"10010101", B"10010101", B"10010101", B"10010101", B"10010101", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010101", B"10010101", B"10010101", B"10010110", B"10010110", B"10010101", B"10010101", B"10010101", B"10010101", B"10010101", B"10010100", B"10010100", B"10010100", B"10010100", B"10010010", B"10010001", B"10001111", B"10010001", B"10001100", B"10001111", B"10010010", B"10001110", B"10000101", B"01110101", B"01100101", B"01011010", B"01011110", B"01110001", B"10001010", B"10010011", B"10001010", B"01111110", B"01111000", B"01111010", B"01111001", B"01111000", B"01111000", B"01110111", B"01110110", B"01110101", B"01110010", B"01110001", B"01101111", B"01101011", B"01101000", B"01100100", B"01100000", B"01011100", B"01011010", B"01011010", B"01010100", B"01000111", B"00110110", B"00111001", B"01000111", B"01001001", B"01001010", B"01001101", B"01001101", B"01110001", B"10001100", B"10001101", B"10001001", B"10001100", B"10001101", B"10001000", B"10000001", B"01111010", B"01110011", B"01011110", B"01011010", B"01001101", B"00110001", B"00100000", B"00010100", B"00011110", B"00011101", B"00010111", B"00010110", B"00010110", B"00110010", B"01001101", B"01101111", B"01101001", B"01100111", B"01100100", B"01100001", B"01100100", B"01110101", B"10001000", B"10001110", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001000", B"10000111", B"10000111", B"10000111", B"10000111", B"10001010", B"10001101", B"10001101", B"10001011", B"10001000", B"10000111", B"10000111", B"10000111", B"10000101", B"10000011", 
B"10000011", B"10000110", B"10001000", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001011", B"10001100", B"10001010", B"01111101", B"01100100", B"01100110", B"01111110", B"10001101", B"10001010", B"10000111", B"10000110", B"10000111", B"10001010", B"10001100", B"10001100", B"10001010", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001010", B"10001100", B"10000011", B"01101011", B"01011011", B"01101001", B"10000011", B"01110101", B"01110010", B"01110000", B"01110001", B"01110000", B"01101111", B"01110000", B"01110000", B"01101000", B"01011110", B"01100100", B"01110101", B"10000000", B"01111110", B"01111001", B"01111000", B"01111000", B"01111001", B"01111001", B"01111010", B"01111010", B"01111010", B"01111010", B"01111010", B"01111010", B"01111010", B"01111001", B"01111001", B"01111001", B"01110110", B"01110101", B"01110110", B"01101111", B"01101011", B"01101001", B"01100101", B"01100101", B"01101000", B"01101011", B"01101100", B"01101100", B"01101110", B"01101011", B"01101001", B"01101000", B"01101000", B"01100101", B"01100011", B"10001011", 
B"10010100", B"10100001", B"10101000", B"10101000", B"10100001", B"10011000", B"10010010", B"10010001", B"10001101", B"10001100", B"10001101", B"10001101", B"10001100", B"10001011", B"10001101", B"10010000", B"10010000", B"10001100", B"10001110", B"10010111", B"10100000", B"10101000", B"10110100", B"10111001", B"10111000", B"11000010", B"11000100", B"10110000", B"10010010", B"10000011", B"10000101", B"10000100", B"10000010", B"01111111", B"01111101", B"01111001", B"01111000", B"01110110", B"01110101", B"01110110", B"01111001", B"01111010", B"01111001", B"01111001", B"01111100", B"01111100", B"01111100", B"01111101", B"01111101", B"01111100", B"01111011", B"01111010", B"01111010", B"01111001", B"01111001", B"01111001", B"01111001", B"01111001", B"01111001", B"01111000", B"01110111", B"01110101", B"01110101", B"01110100", B"01110100", B"01110011", B"01110001", B"01110001", B"01110000", B"01101110", B"01101110", B"01101110", B"01101101", B"01101101", B"01101101", B"01101100", B"01101011", B"01101011", B"01101010", B"01101010", B"01101011", B"01101101", B"01101011", B"01101110", B"01011101", B"00111010", B"01001001", B"01101011", B"01101110", B"01101100", B"01101100", B"01101010", B"01101110", B"01110011", B"01110100", B"01101011", B"01101010", B"01101011", B"01101010", B"01101011", B"01101100", B"01101100", B"01110011", B"01100110", B"01000100", B"00110001", B"00101111", B"00110111", B"00111111", B"01000000", B"01000010", B"00111111", B"00111110", B"00111100", B"00111100", B"00111011", B"00111011", B"00111011", B"00111011", B"00111001", B"00111011", B"00111000", B"00110010", B"00101010", B"00100011", B"00100010", B"00100010", B"00100010", B"00100010", B"00100011", B"00100011", B"00100011", B"00100011", B"00100010", B"00100000", B"00100111", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", 
B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", 
B"01101001", B"01101001", B"01101000", B"01101000", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100100", B"01100101", B"01100101", B"01100101", B"01100111", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101000", B"01101000", B"01100111", B"01100111", B"01101001", B"01101000", B"01100000", B"01011001", B"01100000", B"01101010", B"01100100", B"01101001", B"01101110", B"01101011", B"01100101", B"01100100", B"01101010", B"01110101", B"10000001", B"10010001", B"10011010", B"10100000", B"10100001", B"10011011", B"10010101", B"10010100", B"10010011", B"10010101", B"10010101", B"10010110", B"10011000", B"10011001", B"10011010", B"10011010", B"10011011", B"10011011", B"10011011", B"10011010", B"10011010", B"10011011", B"10011010", B"10011001", B"10010110", B"10010101", B"10010100", B"10010100", B"10010100", B"10010100", B"10010101", B"10010101", B"10010101", B"10010101", B"10010101", B"10010101", B"10010100", B"10010100", B"10010011", B"10010010", B"10010010", B"10010011", B"10010100", B"10010100", B"10010010", B"10010001", B"10010011", B"10010101", B"10010101", B"10010010", B"10001011", B"01111100", B"01101011", B"01011101", B"01010111", B"01011010", B"01110010", B"10000100", B"10001100", B"10001011", B"10000101", B"01111101", B"01111100", B"10000100", B"10001111", B"10001110", B"10001101", B"10001011", B"10001010", B"10000111", B"10000111", B"10001000", B"10000111", B"10000110", B"10000011", B"01111110", B"01111000", B"01110011", B"01110000", B"01110000", B"01100101", B"01001001", B"00100111", B"00100001", B"00101110", B"00111001", B"01000001", B"01001000", B"01001110", B"01101001", B"01110110", B"01110001", B"01101010", B"01101010", B"01101110", B"01101011", B"01001011", B"01000111", B"01001111", B"01001100", B"01010011", B"01010010", B"00111010", B"00100000", B"00011011", B"00110001", B"00101100", B"00100011", B"00101011", B"00110000", B"01000000", B"01010001", B"10000110", B"10000110", B"01111000", B"01101011", B"01100101", B"01100100", B"01110010", B"10000110", B"10001110", B"10001010", B"10001010", B"10001010", B"10001010", B"10001010", B"10001000", B"10000111", B"10000111", B"10000111", B"10000111", B"10001010", B"10001010", B"10001010", B"10000111", B"10000111", B"10000111", B"10000111", B"10000110", B"10000011", B"01111111", 
B"01111111", B"10000011", B"10000110", B"10001010", B"10001011", B"10001100", B"10001100", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001010", B"10001010", B"10001010", B"10001010", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001100", B"10001101", B"10001010", B"01111100", B"01100011", B"01100100", B"01111101", B"10001101", B"10001010", B"10000111", B"10000110", B"10000111", B"10001010", B"10001100", B"10001100", B"10001010", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001010", B"10001100", B"10000011", B"01101011", B"01011011", B"01101001", B"10000011", B"01110011", B"01110001", B"01110000", B"01110000", B"01110000", B"01101111", B"01110000", B"01110000", B"01101000", B"01011110", B"01100011", B"01110101", B"01111111", B"01111101", B"01111000", B"01110111", B"01110111", B"01111000", B"01111000", B"01111001", B"01111001", B"01111010", B"01111001", B"01111001", B"01111001", B"01111000", B"01110111", B"01110111", B"01110110", B"01110011", B"01110001", B"01110010", B"01101110", B"01110000", B"01101110", B"01101010", B"01101010", B"01101100", B"01101110", B"01101100", B"01101100", B"01101100", B"01101010", B"01101001", B"01101000", B"01100111", B"01100101", B"01100101", B"10100111", 
B"10101001", B"10101010", B"10100110", B"10011100", B"10010100", B"10010001", B"10010000", B"10001110", B"10001110", B"10010000", B"10001110", B"10001100", B"10001011", B"10001010", B"10001011", B"10001011", B"10001011", B"10001110", B"10010111", B"10100000", B"10101001", B"10110101", B"10111011", B"10101111", B"10101001", B"10110101", B"10111110", B"10101110", B"10001110", B"01111110", B"10000100", B"10000000", B"01111111", B"01111101", B"01111011", B"01111001", B"01110111", B"01110110", B"01110101", B"01110111", B"01111000", B"01110111", B"01110101", B"01110110", B"01111010", B"01111101", B"01111101", B"01111101", B"01111101", B"01111100", B"01111011", B"01111010", B"01111001", B"01111001", B"01111001", B"01111001", B"01111010", B"01111001", B"01111001", B"01111000", B"01110111", B"01110101", B"01110100", B"01110011", B"01110011", B"01110010", B"01110001", B"01110000", B"01110000", B"01101110", B"01101110", B"01101101", B"01101100", B"01101100", B"01101100", B"01101011", B"01101011", B"01101010", B"01101010", B"01101011", B"01101101", B"01101101", B"01101011", B"01101100", B"01010100", B"00110100", B"01001100", B"01101101", B"01101101", B"01101100", B"01110010", B"01110000", B"01110001", B"01110011", B"01110001", B"01101100", B"01100110", B"01101001", B"01100110", B"01101001", B"01100111", B"01100101", B"01101110", B"01011011", B"00110100", B"00101110", B"00110001", B"00110101", B"00111110", B"00111111", B"01000100", B"00111111", B"00111110", B"00111100", B"00111100", B"00111011", B"00111011", B"00111001", B"00111001", B"00111001", B"00111000", B"00110110", B"00110000", B"00101001", B"00100100", B"00100010", B"00100010", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100010", B"00100000", B"00100111", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", 
B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", 
B"01101010", B"01101001", B"01101001", B"01101000", B"01100111", B"01100111", B"01100101", B"01100101", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01101000", B"01101000", B"01101000", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100101", B"01101000", B"01101000", B"01100000", B"01011001", B"01100000", B"01101111", B"10001010", B"10000111", B"10000101", B"01111111", B"01110111", B"01110000", B"01101010", B"01101001", B"01101011", B"01110101", B"10000001", B"10001110", B"10011000", B"10011000", B"10010101", B"10010011", B"10010010", B"10010100", B"10010100", B"10010101", B"10010110", B"10011000", B"10011001", B"10011010", B"10011011", B"10011011", B"10011100", B"10011101", B"10011101", B"10011101", B"10011100", B"10011010", B"10011000", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010101", B"10010101", B"10010101", B"10010101", B"10010100", B"10010011", B"10010010", B"10001111", B"10001110", B"10001111", B"10010001", B"10010101", B"10010101", B"10010100", B"10010110", B"10010011", B"10001110", B"10001111", B"10000100", B"01110101", B"01100011", B"01010110", B"01011011", B"01101001", B"01110111", B"10000101", B"10001011", B"10001000", B"10000111", B"10000001", B"01111100", B"10000000", B"10001010", B"10001101", B"10001101", B"10001100", B"10001100", B"10001011", B"10001010", B"10001011", B"10001011", B"10001111", B"10010001", B"10010001", B"10001111", B"10001110", B"10001101", B"10001110", B"10001101", B"10001100", B"01110101", B"01001010", B"00101010", B"00100001", B"00100100", B"00100011", B"00101100", B"00110000", B"01001101", B"01010000", B"01000111", B"01000000", B"01000100", B"01001100", B"01010001", B"01010101", B"01011100", B"01110010", B"01111001", B"01111111", B"10000011", B"01100100", B"00111000", B"00101000", B"00111101", B"00111100", B"00110101", B"01000001", B"01000001", B"01000111", B"01010011", B"10001101", B"10001101", B"01111110", B"01110101", B"01101110", B"01100100", B"01110000", B"10001110", B"10001110", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001011", B"10001010", B"10001010", B"10001011", B"10001100", B"10001010", B"10000111", B"10000101", B"10000101", B"10000111", B"10001000", B"10000111", B"10000101", B"10000000", 
B"01111110", B"01111111", B"10000100", B"10001001", B"10001010", B"10001011", B"10001011", B"10001011", B"10001011", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001100", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001110", B"10010000", B"10001010", B"01111100", B"01100011", B"01100100", B"01111101", B"10001100", B"10001001", B"10000110", B"10000110", B"10000111", B"10001010", B"10001100", B"10001100", B"10001010", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001010", B"10001100", B"10000011", B"01101011", B"01011011", B"01101001", B"10000011", B"01110011", B"01110001", B"01110000", B"01110000", B"01110000", B"01101110", B"01110000", B"01110000", B"01101000", B"01011110", B"01100011", B"01110011", B"01111110", B"01111100", B"01110111", B"01110110", B"01110111", B"01110111", B"01111000", B"01111000", B"01111000", B"01111001", B"01111001", B"01111001", B"01111000", B"01111000", B"01110110", B"01110110", B"01110101", B"01110010", B"01110000", B"01110000", B"01110001", B"01110011", B"01110011", B"01110000", B"01110000", B"01110001", B"01101111", B"01101011", B"01101010", B"01101001", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01101001", B"10111100", 
B"10110001", B"10100010", B"10011010", B"10010111", B"10010100", B"10001110", B"10001100", B"10001100", B"10001110", B"10001110", B"10001110", B"10001100", B"10001100", B"10001011", B"10001001", B"10001001", B"10001101", B"10010111", B"10100000", B"10101001", B"10110100", B"10111001", B"10110111", B"10100001", B"10011011", B"10101010", B"10111001", B"10101010", B"10001010", B"01111011", B"10000011", B"01111101", B"01111011", B"01111001", B"01111001", B"01111000", B"01111000", B"01110111", B"01110110", B"01111000", B"01111010", B"01110110", B"01110001", B"01110010", B"01111001", B"01111110", B"01111101", B"01111011", B"01111011", B"01111011", B"01111010", B"01111001", B"01111001", B"01111001", B"01111001", B"01111001", B"01111010", B"01111001", B"01111001", B"01111000", B"01110101", B"01110100", B"01110100", B"01110100", B"01110011", B"01110010", B"01110000", B"01101110", B"01101101", B"01101101", B"01101100", B"01101100", B"01101100", B"01101100", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101100", B"01101110", B"01101110", B"01101101", B"01101100", B"01001100", B"00110000", B"01001110", B"01110001", B"01101101", B"01101110", B"01110111", B"01110010", B"01110010", B"01110011", B"01101101", B"01101011", B"01100011", B"01100110", B"01100101", B"01100111", B"01100111", B"01100101", B"01101101", B"01010011", B"00101001", B"00101010", B"00110001", B"00110010", B"00111001", B"00111011", B"00111111", B"00111100", B"00111011", B"00111001", B"00111000", B"00111000", B"00111000", B"00111000", B"00111000", B"00110111", B"00110110", B"00110010", B"00101110", B"00101001", B"00100100", B"00100011", B"00100010", B"00100010", B"00100010", B"00100011", B"00100011", B"00100011", B"00100011", B"00100010", B"00100000", B"00100111", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", 
B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101100", B"01101100", B"01101100", B"01101011", 
B"01101011", B"01101010", B"01101001", B"01101001", B"01101000", B"01100111", B"01100101", B"01100101", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100101", B"01101000", B"01100111", B"01100000", B"01011001", B"01100000", B"01101111", B"10010010", B"10010001", B"10001110", B"10001101", B"10001011", B"10000111", B"10000000", B"01111000", B"01101111", B"01100111", B"01101010", B"01110010", B"01111010", B"10000001", B"10000101", B"10000110", B"10001000", B"10001000", B"10001000", B"10001000", B"10001010", B"10001010", B"10001100", B"10001101", B"10001111", B"10010010", B"10010101", B"10010110", B"10011000", B"10011001", B"10011001", B"10011000", B"10010110", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010101", B"10010110", B"10010101", B"10010101", B"10010100", B"10010010", B"10010001", B"10001101", B"10001100", B"10001100", B"10001111", B"10010110", B"10011011", B"10011001", B"10010001", B"10000110", B"01111100", B"01110110", B"01101010", B"01100000", B"01011100", B"01011110", B"01101011", B"01111100", B"10001100", B"10001111", B"10001010", B"10000111", B"10000110", B"10000000", B"01111101", B"10000001", B"10001000", B"10001011", B"10001010", B"10001010", B"10001010", B"10001011", B"10001011", B"10001011", B"10001100", B"10001101", B"10001101", B"10001101", B"10001100", B"10001011", B"10001011", B"10001011", B"10001011", B"10001111", B"10001101", B"01100001", B"00111001", B"00110100", B"00101111", B"00100011", B"00110001", B"01100001", B"01110110", B"01110110", B"01110010", B"01110000", B"01110110", B"10000001", B"10001000", B"10001000", B"10001000", B"10010011", B"10010001", B"10001110", B"10010100", B"01111111", B"01001011", B"00101110", B"00111000", B"00110110", B"00101100", B"00110010", B"00110001", B"01000101", B"01100100", B"10001100", B"10001100", B"10000110", B"01111111", B"01110011", B"01011101", B"01100100", B"10001100", B"10001111", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001100", B"10001010", B"10000110", B"10000100", B"10000101", B"10000111", B"10001011", B"10001010", B"10000111", B"10000011", 
B"10000000", B"10000001", B"10000110", B"10001001", B"10001010", B"10001011", B"10001011", B"10001100", B"10001100", B"10001101", B"10001101", B"10001110", B"10001110", B"10010000", B"10010001", B"10010001", B"10010001", B"10010010", B"10010010", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010001", B"10010010", B"10010011", B"10001011", B"01111101", B"01100100", B"01100100", B"01111101", B"10001100", B"10001001", B"10000110", B"10000110", B"10000111", B"10001010", B"10001100", B"10001100", B"10001010", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001010", B"10001100", B"10000011", B"01101011", B"01011011", B"01101001", B"10000011", B"01110011", B"01110001", B"01110000", B"01110000", B"01110000", B"01101111", B"01110000", B"01110000", B"01101000", B"01011110", B"01100010", B"01110010", B"01111101", B"01111100", B"01110111", B"01110110", B"01110111", B"01110111", B"01111000", B"01111000", B"01111000", B"01111001", B"01111010", B"01111001", B"01111001", B"01111000", B"01110110", B"01110110", B"01110101", B"01110001", B"01110000", B"01110000", B"01110000", B"01110010", B"01110010", B"01110000", B"01101111", B"01110000", B"01101110", B"01101010", B"01101001", B"01101000", B"01100101", B"01100101", B"01100100", B"01100011", B"01100111", B"01101010", B"10111000", 
B"10101010", B"10011010", B"10010011", B"10010011", B"10010100", B"10010000", B"10001100", B"10001100", B"10001101", B"10001110", B"10001101", B"10001101", B"10001100", B"10001100", B"10001010", B"10001101", B"10010111", B"10100001", B"10101010", B"10110010", B"10110110", B"10110001", B"10100111", B"10011001", B"10010101", B"10100111", B"10111000", B"10101010", B"10000110", B"01111001", B"10000010", B"01110111", B"01110111", B"01110111", B"01110111", B"01111000", B"01111000", B"01111000", B"01111001", B"01111010", B"01111101", B"01110111", B"01101110", B"01101110", B"01110111", B"01111101", B"01111100", B"01111011", B"01111010", B"01111010", B"01111010", B"01111001", B"01111001", B"01111001", B"01111010", B"01111010", B"01111010", B"01111001", B"01111000", B"01110111", B"01110101", B"01110100", B"01110011", B"01110011", B"01110011", B"01110010", B"01110001", B"01110000", B"01101101", B"01101100", B"01101100", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101110", B"01110010", B"01110011", B"01101001", B"01000010", B"00101100", B"01010001", B"01110101", B"01110010", B"01110000", B"01110111", B"01110010", B"01110001", B"01110011", B"01101101", B"01101010", B"01100010", B"01100101", B"01100101", B"01100111", B"01101010", B"01101010", B"01101011", B"01001011", B"00100101", B"00101001", B"00110000", B"00110000", B"00110001", B"00110010", B"00110111", B"00111001", B"00111000", B"00110111", B"00110111", B"00110111", B"00110111", B"00110111", B"00111000", B"00110110", B"00110100", B"00110000", B"00101101", B"00101001", B"00100110", B"00100010", B"00100001", B"00100010", B"00100011", B"00100011", B"00100011", B"00100011", B"00100011", B"00100010", B"00100000", B"00100111", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", 
B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101100", B"01101100", B"01101100", B"01101100", B"01101100", 
B"01101011", B"01101011", B"01101010", B"01101001", B"01101000", B"01100111", B"01100111", B"01100101", B"01100100", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100101", B"01101000", B"01101000", B"01011110", B"01010110", B"01100001", B"01110000", B"01111110", B"10000100", B"10001100", B"10001110", B"10001110", B"10001101", B"10001101", B"10001100", B"10000001", B"01110110", B"01101110", B"01101010", B"01101000", B"01101111", B"01110001", B"01110111", B"01111001", B"01110111", B"01110111", B"01110111", B"01110110", B"01110110", B"01110110", B"01110110", B"01110111", B"01111010", B"01111110", B"10000000", B"10000011", B"10000101", B"10000110", B"10001011", B"10001110", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010101", B"10010101", B"10010101", B"10010101", B"10010011", B"10010001", B"10001110", B"10001100", B"10001010", B"10001000", B"10010010", B"10011111", B"10011100", B"10010001", B"01111111", B"01110010", B"01101010", B"01100000", B"01100001", B"01100010", B"01101010", B"01110010", B"10000000", B"10001010", B"10010001", B"10001111", B"10001010", B"10000111", B"10000110", B"10000001", B"01111101", B"01111111", B"10000101", B"10000111", B"10000110", B"10000101", B"10000101", B"10000101", B"10000100", B"10000101", B"10000110", B"10010001", B"10010001", B"10001111", B"10001101", B"10001011", B"10000111", B"10000111", B"10000110", B"10001010", B"10001000", B"01011010", B"00110110", B"01000010", B"01000010", B"01000000", B"01001001", B"01111001", B"10000010", B"10000110", B"10001001", B"10001001", B"10001010", B"10001111", B"10010101", B"10001111", B"10000100", B"10001010", B"10001010", B"10000110", B"10000101", B"01110001", B"01000100", B"00101011", B"00110110", B"00110101", B"00101100", B"00101011", B"00101000", B"00111101", B"01100010", B"10000100", B"10001011", B"10001000", B"10000100", B"01110111", B"01011010", B"01100000", B"10000110", B"10010001", B"10001111", B"10001111", B"10001111", B"10001111", B"10001111", B"10001110", B"10001110", B"10001101", B"10001100", B"10001100", B"10001011", B"10000111", B"10000100", B"10000011", B"10000100", B"10000111", B"10001010", B"10001011", B"10001010", B"10000111", 
B"10000111", B"10001000", B"10001100", B"10001101", B"10001101", B"10001110", B"10001110", B"10010000", B"10010000", B"10010000", B"10010001", B"10010001", B"10010010", B"10010010", B"10010010", B"10010011", B"10010011", B"10010011", B"10010011", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010011", B"10001011", B"01111011", B"01100010", B"01100011", B"01111100", B"10001011", B"10001001", B"10000110", B"10000101", B"10000111", B"10001010", B"10001100", B"10001100", B"10001010", B"10001001", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001011", B"10000010", B"01101010", B"01011010", B"01101000", B"10000010", B"01110011", B"01110001", B"01110000", B"01110001", B"01110000", B"01101111", B"01110000", B"01110000", B"01101000", B"01011110", B"01100001", B"01110001", B"01111100", B"01111010", B"01110111", B"01110110", B"01110111", B"01110111", B"01111000", B"01111000", B"01111001", B"01111010", B"01111010", B"01111010", B"01111001", B"01111000", B"01110110", B"01110101", B"01110011", B"01110001", B"01110000", B"01101111", B"01101110", B"01101011", B"01101011", B"01101001", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100101", B"01100100", B"01100011", B"01100011", B"01100111", B"01101100", B"10100111", 
B"10100001", B"10011001", B"10010100", B"10010001", B"10010001", B"10001110", B"10001101", B"10001100", B"10001101", B"10001110", B"10001101", B"10001100", B"10001101", B"10010000", B"10010001", B"10011000", B"10100011", B"10101101", B"10110101", B"10110110", B"10110000", B"10100101", B"10010111", B"10010101", B"10010100", B"10101010", B"10111100", B"10101010", B"10000100", B"01111000", B"01111111", B"01110100", B"01110101", B"01110101", B"01110110", B"01110111", B"01111000", B"01111001", B"01111100", B"01111110", B"01111110", B"01111000", B"01110000", B"01110000", B"01110111", B"01111100", B"01111010", B"01111011", B"01111001", B"01111010", B"01111010", B"01111010", B"01111011", B"01111011", B"01111011", B"01111010", B"01111010", B"01111001", B"01111000", B"01110111", B"01110100", B"01110100", B"01110011", B"01110011", B"01110011", B"01110010", B"01110001", B"01110000", B"01101110", B"01101101", B"01101100", B"01101011", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101010", B"01101110", B"01110011", B"01111000", B"01100110", B"00111011", B"00101100", B"01010111", B"01111011", B"01110111", B"01110010", B"01110101", B"01110001", B"01110000", B"01110010", B"01101110", B"01101101", B"01100110", B"01100111", B"01101010", B"01101010", B"01101011", B"01101110", B"01100101", B"01000010", B"00100100", B"00100111", B"00101111", B"00101110", B"00101110", B"00110000", B"00110100", B"00110101", B"00110101", B"00110101", B"00110101", B"00110110", B"00110110", B"00110110", B"00110111", B"00110110", B"00110010", B"00101111", B"00101011", B"00101001", B"00100110", B"00100011", B"00100001", B"00100000", B"00100001", B"00100010", B"00100010", B"00100010", B"00100010", B"00100001", B"00011111", B"00100111", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", 
B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101100", B"01101100", B"01101100", B"01101100", B"01101100", 
B"01101011", B"01101011", B"01101010", B"01101001", B"01101000", B"01100111", B"01100101", B"01100101", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100101", B"01101000", B"01101001", B"01011110", B"01010101", B"01100001", B"01110001", B"01111111", B"10001011", B"10010110", B"10010100", B"10001100", B"10000110", B"10000111", B"10001100", B"10001101", B"10000111", B"01111111", B"01111001", B"01111001", B"01111000", B"01110011", B"01110011", B"01110010", B"01110001", B"01110001", B"01110000", B"01101111", B"01101110", B"01101100", B"01101011", B"01101011", B"01101011", B"01101011", B"01101010", B"01101010", B"01101011", B"01101100", B"01110010", B"10001000", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010100", B"10010101", B"10010101", B"10010101", B"10010101", B"10010011", B"10010001", B"10001110", B"10001011", B"10001000", B"10001011", B"10010011", B"10011010", B"10001111", B"01111101", B"01101001", B"01100100", B"01101100", B"01011110", B"01100100", B"01110000", B"10000000", B"10001101", B"10010010", B"10001110", B"10001011", B"10001010", B"10001000", B"10000110", B"10000111", B"10000100", B"01111101", B"01111110", B"10000110", B"10001010", B"10001000", B"10000111", B"10000110", B"10000110", B"10000110", B"10000110", B"10000111", B"10001000", B"10001010", B"10001010", B"10001010", B"10001000", B"10000111", B"10001000", B"10000111", B"10010100", B"10010001", B"01100011", B"00111001", B"00111011", B"00111100", B"00111010", B"01000000", B"01110111", B"10000100", B"10001100", B"10010010", B"10010000", B"10001010", B"10000111", B"10001000", B"10001010", B"01111110", B"10000111", B"10010011", B"10001100", B"01110110", B"01010110", B"00111001", B"00110011", B"00111111", B"00111111", B"00111100", B"00111110", B"00111100", B"01000100", B"01011010", B"01111100", B"10000111", B"10000101", B"10000001", B"01111010", B"01100011", B"01100111", B"10000110", B"10010011", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010010", B"10010011", B"10010011", B"10010011", B"10010001", B"10001101", B"10001011", B"10001010", B"10001011", B"10001101", B"10001111", B"10010001", B"10010001", B"10010001", 
B"10010010", B"10010011", B"10010100", B"10010010", B"10010001", B"10010001", B"10010000", B"10010000", B"10010000", B"10010000", B"10010000", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001101", B"10001101", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10001110", B"10010000", B"10010001", B"10001001", B"01111000", B"01100000", B"01100001", B"01111001", B"10001010", B"10001010", B"10000110", B"10000101", B"10000111", B"10001010", B"10001100", B"10001100", B"10001010", B"10001001", B"10001001", B"10001001", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000110", B"10000110", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001010", B"10000000", B"01101001", B"01011010", B"01100111", B"10000000", B"01110010", B"01110001", B"01110000", B"01110001", B"01110000", B"01101111", B"01110000", B"01110000", B"01101000", B"01011101", B"01100001", B"01101111", B"01111001", B"01111001", B"01110111", B"01110110", B"01110111", B"01110111", B"01111000", B"01111000", B"01111000", B"01111010", B"01111010", B"01111010", B"01111001", B"01110111", B"01110101", B"01110101", B"01110011", B"01110000", B"01101111", B"01101111", B"01101011", B"01100111", B"01100100", B"01100101", B"01100011", B"01100000", B"01100000", B"01100011", B"01100100", B"01100101", B"01100111", B"01100111", B"01100101", B"01100101", B"01101011", B"01110001", B"10100000", 
B"10011001", B"10010011", B"10010001", B"10001110", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10001101", B"10010000", B"10010101", B"10011111", B"10101000", B"10101111", B"10110101", B"10110111", B"10110010", B"10100111", B"10011000", B"10001100", B"10010001", B"10010000", B"10110100", B"11000000", B"10101011", B"01111111", B"01111100", B"01111100", B"01110101", B"01110010", B"01110101", B"01110110", B"01110111", B"01111001", B"01111100", B"01111111", B"10000000", B"10000000", B"01111010", B"01110011", B"01110011", B"01111000", B"01111110", B"01111111", B"01111110", B"01111010", B"01111011", B"01111100", B"01111100", B"01111110", B"01111100", B"01111100", B"01111011", B"01111010", B"01111001", B"01110111", B"01110101", B"01110100", B"01110011", B"01110011", B"01110011", B"01110011", B"01110010", B"01110001", B"01101110", B"01101101", B"01101100", B"01101011", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101101", B"01110011", B"01111001", B"01100010", B"00111000", B"00110011", B"01011111", B"01111110", B"01111010", B"01110010", B"01110011", B"01110000", B"01101110", B"01110001", B"01110010", B"01101111", B"01101011", B"01101011", B"01101110", B"01101011", B"01101011", B"01101111", B"01011010", B"00110110", B"00100100", B"00100101", B"00101101", B"00101110", B"00101011", B"00110000", B"00110010", B"00110101", B"00110100", B"00110100", B"00110100", B"00110100", B"00110100", B"00110100", B"00110101", B"00110101", B"00110001", B"00101110", B"00101010", B"00100111", B"00100011", B"00100001", B"00100000", B"00100000", B"00100000", B"00100001", B"00100001", B"00100001", B"00100001", B"00100000", B"00011101", B"00100110", B"01000010", B"01011111", B"01100110", B"01100011", B"01100010", B"01100010", B"01100010", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100000", B"01100001", B"01100001", B"01100010", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100100", B"01100011", B"01100011", 
B"01100011", B"01100011", B"01100011", B"01100010", B"01100010", B"01100010", B"01100011", B"01100011", B"01100011", B"01100011", B"01100100", B"01100100", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100101", B"01100100", B"01100100", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100101", B"01100101", B"01100101", B"01100101", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101001", B"01101001", B"01101001", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101010", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", B"01101011", 
B"01101011", B"01101010", B"01101010", B"01101001", B"01101000", B"01100111", B"01100101", B"01100101", B"01100100", B"01100100", B"01100100", B"01100101", B"01100101", B"01100111", B"01100111", B"01101000", B"01101000", B"01101000", B"01101000", B"01101000", B"01100111", B"01101000", B"01101001", B"01100111", B"01100100", B"01101000", B"01101001", B"01011101", B"01010100", B"01100011", B"10000100", B"10010100", B"10011000", B"10011000", B"10010101", B"10010001", B"10001101", B"10001011", B"10001011", B"10001101", B"10001111", B"10001110", B"10001100", B"10001010", B"10000110", B"10000100", B"10000110", B"10000111", B"10001000", B"10001010", B"10001011", B"10001011", B"10000110", B"01111101", B"01110110", B"01101001", B"01101001", B"01101000", B"01101001", B"01101000", B"01100111", B"01100100", B"01100011", B"01101000", B"01110101", B"10001010", B"10001110", B"10010100", B"10011000", B"10010110", B"10010101", B"10010100", B"10010100", B"10010100", B"10010011", B"10010011", B"10010010", B"10010001", B"10010001", B"10001111", B"10010010", B"10000101", B"01101001", B"01011101", B"01100011", B"01110001", B"01110011", B"01111010", B"10000101", B"10001110", B"10010001", B"10010010", B"10010010", B"10001111", B"10001101", B"10001010", B"10000111", B"10000101", B"10001000", B"10000100", B"01111101", B"01111111", B"10000110", B"10001010", B"10001000", B"10001000", B"10000111", B"10000110", B"10000110", B"10000111", B"10001010", B"10001010", B"10000111", B"10000101", B"10001010", B"10001111", B"10010011", B"10010010", B"10001011", B"10010101", B"10000000", B"01010000", B"00111011", B"01000100", B"00110011", B"00101110", B"01001110", B"10000011", B"10001100", B"10010000", B"10001110", B"10001011", B"10000111", B"10001000", B"10001000", B"10001111", B"10001000", B"10001101", B"10010001", B"01111001", B"01010100", B"00111000", B"00110001", B"00111100", B"01001000", B"01001111", B"01010110", B"01011101", B"01011101", B"01011100", B"01100100", B"01110011", B"01111110", B"10000101", B"10000111", B"10000000", B"01101010", B"01100000", B"01101000", B"01111010", B"01111111", B"10000101", B"10001010", B"10001101", B"10001111", B"10010001", B"10010010", B"10010011", B"10010001", B"10001110", B"10001011", B"10000110", B"10000001", B"01111111", B"01111111", B"01111111", B"01111111", B"01111110", B"01111110", B"01111101", 
B"01111100", B"01111100", B"01111010", B"01111000", B"01111001", B"01111011", B"01111011", B"01111011", B"01111011", B"01111011", B"01111001", B"01111001", B"01111001", B"01111001", B"01111001", B"01111000", B"01111000", B"01111000", B"01111000", B"01111000", B"01111000", B"01111000", B"01111000", B"01111000", B"01111000", B"01111000", B"01111001", B"01111011", B"01111111", B"10000010", B"10000100", B"10000110", B"10001001", B"10001010", B"10001001", B"01111111", B"01101110", B"01011010", B"01011111", B"01110010", B"10000111", B"10001010", B"10000110", B"10000110", B"10000111", B"10001010", B"10001011", B"10001011", B"10001010", B"10001010", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000110", B"10000110", B"10000110", B"10000110", B"10000110", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10001001", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000111", B"10000110", B"10000101", B"10000111", B"01111111", B"01101000", B"01011011", B"01100100", B"01101111", B"01110000", B"01101111", B"01101111", B"01110000", B"01101111", B"01101110", B"01101111", B"01110000", B"01101000", B"01011100", B"01011110", B"01101110", B"01111000", B"01111000", B"01110110", B"01110110", B"01110111", B"01111000", B"01111000", B"01111000", B"01111001", B"01111010", B"01111010", B"01111010", B"01111001", B"01110111", B"01110101", B"01110011", B"01110010", B"01110000", B"01101111", B"01110000", B"01101010", B"01100011", B"01100011", B"01100111", B"01100011", B"01011100", B"01011100", B"01100001", B"01100011", B"01100100", B"01101000", B"01101010", B"01101001", B"01101010", B"01110001", B"01110110"   );

    constant KERNEL_DATA_WIDTH: positive := 16;
 --   constant KERNEL_ADDR_WIDTH: positive := 10;
    constant KERNEL_SIZE: positive := 9;

    constant IMG_BRAM_SIZE: positive := 2160;

    type rom_type is array(0 to KERNEL_SIZE - 1) of std_logic_vector(KERNEL_DATA_WIDTH - 1 downto 0);
    constant KERNEL_CONTENT: rom_type := (
    B"0000100110011101",
    B"0000111111011010",
    B"0000100110011101",
    B"0000111111011010",
    B"0001101000100011",
    B"0000111111011010",
    B"0000100110011101",
    B"0000111111011010",
    B"0000100110011101"
    );

    signal clk_s, reset_s, start_s, ready_s: std_logic;
    signal X_img_data_s: std_logic_vector(7 downto 0);
    signal X_img_addr_s: std_logic_vector(14 downto 0);
    signal X_img_en_s: std_logic;
    signal X_img_we_s: std_logic_vector(3 downto 0);
    signal kernel_en_s: std_logic;
    signal kernel_we_s: std_logic_vector(3 downto 0);
    signal kernel_addr_s: std_logic_vector(9 downto 0);
    signal kernel_data_s: std_logic_vector(15 downto 0);
    signal kernel_size_in_s: std_logic_vector(4 downto 0);
    signal dram_we_s: std_logic;
    signal dram_data_s: std_logic_vector(7 downto 0);
    signal dram_addr_s : std_logic_vector(21 downto 0);
    signal axi_read_init_s, axi_rready_s, axi_read_last_s, axi_rvalid_s: std_logic;
    signal axi_burst_len_s: std_logic_vector(7 downto 0);
    signal axi_raddr_s: std_logic_vector(21 downto 0);
    signal img_bram_waddr_s: std_logic_vector(14 downto 0);
    signal img_wdata_s: std_logic_vector(7 downto 0);
    signal axi_write_init_s: std_logic;

begin

clk_gen: process
begin
    clk_s <= '0', '1' after 5 ns;
    wait for 10 ns;
end process;

stim_gen: process
begin
    reset_s <= '1';
    start_s <= '0';
    wait for 25 ns;
    reset_s <= '0';
    wait until falling_edge(clk_s);
    X_img_en_s <= '1';
    X_img_we_s <= "1111";
    for j in 0 to 3 loop
    for i in 0 to 720 loop
        X_img_addr_s <= conv_std_logic_vector(j*720+i, X_img_addr_s'length);
        X_img_data_s <= DRAM_CONTENT(j*720 + i);
        wait until falling_edge(clk_s);
    end loop;
    end loop;
    X_img_en_s <= '0';
    X_img_we_s <= "0000";
    
    wait until falling_edge(clk_s);
    kernel_en_s <= '1';
    kernel_we_s <= "1111";
    for i in 0 to KERNEL_SIZE - 1 loop
        kernel_addr_s <= conv_std_logic_vector(i, kernel_addr_s'length);
        kernel_data_s <= KERNEL_CONTENT(i);
        wait until falling_edge(clk_s);
    end loop;
    kernel_en_s <= '0';
    kernel_we_s <= "0000";    

    reset_s <= '1';    
    wait until falling_edge(clk_s);
    reset_s <= '0';
    start_s <= '1';
    axi_read_last_s <= '0';
    axi_rvalid_s <= '0';
    kernel_size_in_s <= "00011";
    wait until falling_edge(clk_s);
    start_s <= '0';
    
    wait until axi_read_init_s = '1';
    wait until rising_edge(clk_s);
    axi_rvalid_s <= '1';
    
    for i in 0 to 255 loop
        img_wdata_s <= DRAM_CONTENT(2160+i);
        if(i = 255) then
            axi_read_last_s <= '1';        
        end if;
        wait until rising_edge(clk_s);   
        
    end loop;

    axi_read_last_s <= '0';
    axi_rvalid_s <= '0';
    
    wait until axi_read_init_s = '1';
    wait until rising_edge(clk_s);
    axi_rvalid_s <= '1';
 
 
    for i in 256 to 511 loop
        img_wdata_s <= DRAM_CONTENT(2160+i);
        if(i = 511) then
            axi_read_last_s <= '1';        
        end if;
        wait until rising_edge(clk_s);   
        
    end loop;

    axi_read_last_s <= '0';
    axi_rvalid_s <= '0';
    
    wait until axi_read_init_s = '1';
    wait until rising_edge(clk_s);
    axi_rvalid_s <= '1';    

    for i in 512 to 719 loop
        img_wdata_s <= DRAM_CONTENT(2160+i);
        if(i = 719) then
            axi_read_last_s <= '1';        
        end if;
        wait until rising_edge(clk_s);   
        
    end loop;


    axi_read_last_s <= '0';
    axi_rvalid_s <= '0';
    
    wait until ready_s = '1';
        
    wait;
end process;


--Ovo je DUV

duv: entity work.apply_gaussian_top 
Port map( 
    ---------- Clocking and reset interface----------
    clk => clk_s,
    reset => reset_s,

    ---------- Input ------------
    kernel_size_i => kernel_size_in_s,

    ---------- Command interface ----------
    start => start_s,

    ---------- IPB to DRAM interface  ----------
   -- dram_we_o => dram_we_s,
    dram_waddr_o => dram_addr_s,
    dram_wdata_o => dram_data_s,

    ---- IMG BRAM to DRAM -----
    img_en_i => X_img_en_s,
    img_we_i => X_img_we_s,
    img_waddr_b_i => X_img_addr_s,
    img_wdata_b_i => X_img_data_s,
    
    ---- IPB READS DRAM ----
    img_wdata_i => img_wdata_s,

    ---- KERNEL BRAM to CPU ----
    kernel_en_i => kernel_en_s,
    kernel_we_i => kernel_we_s,
    kernel_waddr_i => kernel_addr_s,
    kernel_wdata_i => kernel_data_s,

    ---------- Status interface ----------
    ready_o => ready_s, 
    
    -- AXI read dram --
    axi_read_init_o => axi_read_init_s,
    axi_burst_len_o => axi_burst_len_s,
    --axi_rready_o => axi_rready_s,
    axi_read_last_i => axi_read_last_s,
    axi_raddr_o => axi_raddr_s,
    axi_rvalid_i => axi_rvalid_s,
    
    -- AXI writes dram --
    axi_write_init_o => axi_write_init_s
           
  );

end Behavioral;
